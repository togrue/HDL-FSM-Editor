-- Filename: regression2_e.vhd
-- Created by HDL-FSM-Editor
library ieee;
use ieee.std_logic_1164.all;

entity regression2 is
    port (
        res_i : in std_logic;
        clk_i : in std_logic
    );
end entity;
